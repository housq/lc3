`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    05:17:23 03/22/2014 
// Design Name: 
// Module Name:    LC3_FSM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module LC3_FSM(
		input						clk,
		input						reset,
		input						Priv,
		input						BEN,
		input			[15:11]	IR,
		input						R,
		input						INT,
		
		output	reg[39:0]	CONTROL
    );
	 
	wire				[49:0]	SIGNALS		[63:0];	

	reg				[5:0]		CS,NS;
	reg				[5:0]		J;
	reg				[2:0]		COND;
	reg							IRD;
	
assign SIGNALS[0 ] = 50'b00100100100000000000000000000000000000000000000000;
assign SIGNALS[1 ] = 50'b00000100100000110000000010000000000100000000000000;
assign SIGNALS[2 ] = 50'b00000110011000000000000001000000000001000100000000;
assign SIGNALS[3 ] = 50'b00000101111000000000000001000000000001000100000000;
assign SIGNALS[4 ] = 50'b00110101000000100000001000000000010000000000000000;
assign SIGNALS[5 ] = 50'b00000100100000110000000010000000000100000000001000;
assign SIGNALS[6 ] = 50'b00000110011000000000000001000000000110100100000000;
assign SIGNALS[7 ] = 50'b00000101111000000000000001000000000110100100000000;
assign SIGNALS[8 ] = 50'b01001001001000000000000010000000001000000000011000;
assign SIGNALS[9 ] = 50'b00000100100000110000000010000000000100000000010000;
assign SIGNALS[10] = 50'b00000110001000000000000001000000000001000100000000;
assign SIGNALS[11] = 50'b00000111011000000000000001000000000001000100000000;
assign SIGNALS[12] = 50'b00000100100000001000000000000010000110000000000000;
assign SIGNALS[13] = 50'b01001001010100000010010000001000000000000010000000;
assign SIGNALS[14] = 50'b00000100100000110000000001000000000001000100000000;
assign SIGNALS[15] = 50'b00000111001000000000000001000000000000000000000000;
assign SIGNALS[16] = 50'b00010100000000000000000000000000000000000000000110;
assign SIGNALS[17] = 50'b00000000000000000000000000000000000000000000000000;
assign SIGNALS[18] = 50'b01011000011000001000001000000000000000000000000000;
assign SIGNALS[19] = 50'b00000000000000000000000000000000000000000000000000;
assign SIGNALS[20] = 50'b00000100100000101000001000000010010110000000000000;
assign SIGNALS[21] = 50'b00000100100000001000000000000010000001100000000000;
assign SIGNALS[22] = 50'b00000100100000001000000000000010000001000000000000;
assign SIGNALS[23] = 50'b00000100000100000000000010000000000000000000011000;
assign SIGNALS[24] = 50'b00010110000100000000000000000000000000000000000100;
assign SIGNALS[25] = 50'b00010110010100000000000000000000000000000000000100;
assign SIGNALS[26] = 50'b00000110011000000000000100000000000000000000000000;
assign SIGNALS[27] = 50'b00000100100000110000000100000000000000000000000000;
assign SIGNALS[28] = 50'b00010111000100100000001000000000010000000000000100;
assign SIGNALS[29] = 50'b00010111010100000000000000000000000000000000000100;
assign SIGNALS[30] = 50'b00000100100000001000000100000001000000000000000000;
assign SIGNALS[31] = 50'b00000101111000000000000100000000000000000000000000;
assign SIGNALS[32] = 50'b10000000000001000000000000000000000000000000000000;
assign SIGNALS[33] = 50'b00011000010100000000000000000000000000000000000100;
assign SIGNALS[34] = 50'b01001100110000100000000000000100101000000000000000;
assign SIGNALS[35] = 50'b00001000000010000000000100000000000000000000000000;
assign SIGNALS[36] = 50'b00011001000100000000000000000000000000000000000100;
assign SIGNALS[37] = 50'b00001010011000100000000000000100101000001000000000;
assign SIGNALS[38] = 50'b00001001110000001000000100000001000000000000000000;
assign SIGNALS[39] = 50'b00001010001000100000000000000100101000000000000000;
assign SIGNALS[40] = 50'b00011010000100000000000000000000000000000000000100;
assign SIGNALS[41] = 50'b00011010010000000000000000000000000000000000100110;
assign SIGNALS[42] = 50'b00001000100000010110000100000000000000000000000000;
assign SIGNALS[43] = 50'b00001011110100000000000000010000000000000000000000;
assign SIGNALS[44] = 50'b00001011010100000010010000001000000000000001000000;
assign SIGNALS[45] = 50'b00001001010000100000100000000100101000010000000000;
assign SIGNALS[46] = 50'b00000000000000000000000000000000000000000000000000;
assign SIGNALS[47] = 50'b00001100001000100000000000000100101000001000000000;
assign SIGNALS[48] = 50'b00011100000000000000000000000000000000000000000110;
assign SIGNALS[49] = 50'b01001001010100000110010000001000000000000000000000;
assign SIGNALS[50] = 50'b00001101001000000000000000100000000000000000000000;
assign SIGNALS[51] = 50'b00000100100000000000000000000000000000000000000000;
assign SIGNALS[52] = 50'b00011101000100000000000000000000000000000000000100;
assign SIGNALS[53] = 50'b00000000000000000000000000000000000000000000000000;
assign SIGNALS[54] = 50'b00000100100000001000000100000001000000000000000000;
assign SIGNALS[55] = 50'b00000000000000000000000000000000000000000000000000;
assign SIGNALS[56] = 50'b00000000000000000000000000000000000000000000000000;
assign SIGNALS[57] = 50'b00000000000000000000000000000000000000000000000000;
assign SIGNALS[58] = 50'b00000000000000000000000000000000000000000000000000;
assign SIGNALS[59] = 50'b00000100100000100001000000000100101000011000000000;
assign SIGNALS[60] = 50'b00000000000000000000000000000000000000000000000000;
assign SIGNALS[61] = 50'b00000000000000000000000000000000000000000000000000;
assign SIGNALS[62] = 50'b00000000000000000000000000000000000000000000000000;
assign SIGNALS[63] = 50'b00000000000000000000000000000000000000000000000000;
	
	
	always@(*)	begin
		if(reset)
				NS=6'd18;
		else if(IRD)
				NS={2'b00,IR[15:12]};
		else 
				NS=	{J[5],
						 J[4]|( COND[2]& ~COND[1]& COND[0] &INT)		,
						 J[3]|( COND[2]& ~COND[1]&~COND[0] &Priv)	,
						 J[2]|(~COND[2]&  COND[1]&~COND[0] &BEN)		,
						 J[1]|(~COND[2]& ~COND[1]& COND[0] &R)			,
						 J[0]|(~COND[2]&  COND[1]& COND[0] &IR[11])	
						};
						
	end
	
	
	always@(posedge clk)	begin
		CS<=NS;
	end
	
	always@(posedge clk)	begin
			{IRD,COND,J,CONTROL}<=SIGNALS[NS];
	end
	
	

endmodule
